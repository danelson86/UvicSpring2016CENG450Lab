----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    01:26:03 03/01/2016 
-- Design Name: 
-- Module Name:    EXtoMem_pipeline - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity EXtoMem_pipeline is
	Port(
			CLK : in STD_LOGIC:='0';
			RST : in STD_LOGIC:='0'; 
			
			Data1 : in	STD_LOGIC_VECTOR (15 downto 0):= X"0000";
			Data2  : in		STD_LOGIC_VECTOR (15 downto 0):= X"0000";
			WB_rqst_ADDR : in	 STD_LOGIC_VECTOR (2 downto 0):="000";
			microcode :in std_logic_vector(3 downto 0) := "0000";
			
			Data1x : out	STD_LOGIC_VECTOR (15 downto 0):= X"0000";
			Data2x  : out	STD_LOGIC_VECTOR (15 downto 0):= X"0000";
			WB_rqst_ADDRx : out STD_LOGIC_VECTOR (2 downto 0):="000";
			microcodeX : out std_logic_vector(3 downto 0) := "0000");
			
end EXtoMem_pipeline;

architecture Behavioral of EXtoMem_pipeline is

component pipeline_16bit is
		Port(
			clk : in STD_LOGIC:='0';
			rst : in STD_LOGIC:='0';
			input : in STD_LOGIC_VECTOR(15 downto 0):= X"0000";
			output : out STD_LOGIC_VECTOR(15 downto 0):= X"0000");
	end component;
	
	component pipeline_5deep_3bit is
		Port(
			clk : in STD_LOGIC:='0';
			rst : in STD_LOGIC:='0';
			input : in STD_LOGIC_VECTOR(2 downto 0):="000";
			output : out STD_LOGIC_VECTOR(2 downto 0):="000");
	end component;
	
	component pipeline_4bit is
		Port(
			clk : in STD_LOGIC := '0';
			rst : in STD_LOGIC := '0';
			input : in STD_LOGIC_VECTOR(3 downto 0):= X"0";
			output : out STD_LOGIC_VECTOR(3 downto 0):= X"0");
	end component;
	


begin


	data1pipe : pipeline_16bit port map(clk,rst,data1,data1x);
	data2pipe : pipeline_16bit port map(clk,rst,data2,data2x);
	wb_rqst_addr_pipe : pipeline_5deep_3bit port map (clk,rst,WB_Rqst_Addr,WB_Rqst_AddrX);
	microcodePipe : pipeline_4bit port map(clk,rst,microcode,microcodeX);
	
end Behavioral;

